
module FetchModule (input clk, input reset, input [31:0] next_pc_in, output [24:0] bundle_out);



endmodule