
module DecodeModule (input clk, input reset, input bundle_in [24:0], output reg [12:0] bundle_out,
		input [31:0] pc_seq_in, input [31:0] pc_seq_2_in, output [31:0] pc_seq_out);

endmodule