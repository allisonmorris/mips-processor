
module MemoryModule (input clk, input reset, input [6:0] bundle_in, output reg [1:0] bundle_out,
		input [31:0] pc_seq_in, output [31:0] pc_seq_out);

endmodule